module test (
);




endmodule
